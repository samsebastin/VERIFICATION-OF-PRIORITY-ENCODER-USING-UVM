

////////////////////////////////////////////////////////////////////////////////////////////////////

module top;

	import uvm_pkg::*;
	
	import pe_pkg::*;

	pe_vif vif();
	
	pe dut(.in(vif.in),.out(vif.out));

initial
begin
	uvm_config_db#(virtual pe_vif)::set(null,"*","pe_vif",vif);
	run_test("test");
end

endmodule

/////////////////////////////////////////////////////////////////////////////////////////////////