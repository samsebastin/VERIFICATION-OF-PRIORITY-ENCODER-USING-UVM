

//////////////////////////////////////////////////////////////////////////////////////////

interface pe_vif();

	bit [3:0] in;
	bit [1:0] out;
	
	modport WR_DRV_MP(output in);
	modport WR_MON_MP(input in);
	modport RD_MON_MP(input out);
	
endinterface

//////////////////////////////////////////////////////////////////////////////////////////