

//////////////////////////////////////////////////////////////////////////////////////////

class write_config extends uvm_object;

	`uvm_object_utils(write_config)
	
	function new(string name="write_config");
		super.new(name);
	endfunction
	
	virtual pe_vif vif;
	uvm_active_passive_enum is_active;
	
endclass

////////////////////////////////////////////////////////////////////////////////////////